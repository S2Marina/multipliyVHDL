-- MySoc.vhd

-- Generated using ACDS version 13.0sp1 232 at 2022.03.23.11:27:48

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MySoc is
	port (
		clk_clk       : in  std_logic                     := '0';             --   clk.clk
		reset_reset_n : in  std_logic                     := '0';             -- reset.reset_n
		go_export     : out std_logic;                                        --    go.export
		prt_export    : in  std_logic                     := '0';             --   prt.export
		res_export    : in  std_logic_vector(11 downto 0) := (others => '0'); --   res.export
		mult_export   : out std_logic_vector(5 downto 0);                     --  mult.export
		m_export      : out std_logic_vector(5 downto 0)                      --     m.export
	);
end entity MySoc;

architecture rtl of MySoc is
	component MySoc_nios is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(17 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component MySoc_nios;

	component MySoc_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component MySoc_ram;

	component MySoc_jtag is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component MySoc_jtag;

	component MySoc_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component MySoc_sysid;

	component MySoc_m is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(5 downto 0)                      -- export
		);
	end component MySoc_m;

	component MySoc_res is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(11 downto 0) := (others => 'X')  -- export
		);
	end component MySoc_res;

	component MySoc_prt is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component MySoc_prt;

	component MySoc_go is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component MySoc_go;

	component MySoc_performance_counter_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component MySoc_performance_counter_0;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(92 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component altera_merlin_slave_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(17 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(92 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(93 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_agent;

	component altera_avalon_sc_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(93 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component altera_avalon_sc_fifo;

	component MySoc_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(92 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component MySoc_addr_router;

	component MySoc_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(92 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component MySoc_addr_router_001;

	component MySoc_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(92 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component MySoc_id_router;

	component MySoc_id_router_005 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(92 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component MySoc_id_router_005;

	component MySoc_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(92 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(92 downto 0);                    -- data
			src1_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(92 downto 0);                    -- data
			src2_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(92 downto 0);                    -- data
			src3_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic;                                        -- endofpacket
			src4_ready         : in  std_logic                     := 'X';             -- ready
			src4_valid         : out std_logic;                                        -- valid
			src4_data          : out std_logic_vector(92 downto 0);                    -- data
			src4_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src4_startofpacket : out std_logic;                                        -- startofpacket
			src4_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component MySoc_cmd_xbar_demux;

	component MySoc_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(92 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(92 downto 0);                    -- data
			src1_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(92 downto 0);                    -- data
			src2_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(92 downto 0);                    -- data
			src3_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic;                                        -- endofpacket
			src4_ready         : in  std_logic                     := 'X';             -- ready
			src4_valid         : out std_logic;                                        -- valid
			src4_data          : out std_logic_vector(92 downto 0);                    -- data
			src4_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src4_startofpacket : out std_logic;                                        -- startofpacket
			src4_endofpacket   : out std_logic;                                        -- endofpacket
			src5_ready         : in  std_logic                     := 'X';             -- ready
			src5_valid         : out std_logic;                                        -- valid
			src5_data          : out std_logic_vector(92 downto 0);                    -- data
			src5_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src5_startofpacket : out std_logic;                                        -- startofpacket
			src5_endofpacket   : out std_logic;                                        -- endofpacket
			src6_ready         : in  std_logic                     := 'X';             -- ready
			src6_valid         : out std_logic;                                        -- valid
			src6_data          : out std_logic_vector(92 downto 0);                    -- data
			src6_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src6_startofpacket : out std_logic;                                        -- startofpacket
			src6_endofpacket   : out std_logic;                                        -- endofpacket
			src7_ready         : in  std_logic                     := 'X';             -- ready
			src7_valid         : out std_logic;                                        -- valid
			src7_data          : out std_logic_vector(92 downto 0);                    -- data
			src7_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src7_startofpacket : out std_logic;                                        -- startofpacket
			src7_endofpacket   : out std_logic;                                        -- endofpacket
			src8_ready         : in  std_logic                     := 'X';             -- ready
			src8_valid         : out std_logic;                                        -- valid
			src8_data          : out std_logic_vector(92 downto 0);                    -- data
			src8_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src8_startofpacket : out std_logic;                                        -- startofpacket
			src8_endofpacket   : out std_logic;                                        -- endofpacket
			src9_ready         : in  std_logic                     := 'X';             -- ready
			src9_valid         : out std_logic;                                        -- valid
			src9_data          : out std_logic_vector(92 downto 0);                    -- data
			src9_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src9_startofpacket : out std_logic;                                        -- startofpacket
			src9_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component MySoc_cmd_xbar_demux_001;

	component MySoc_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(92 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component MySoc_cmd_xbar_mux;

	component MySoc_rsp_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(92 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(92 downto 0);                    -- data
			src1_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component MySoc_rsp_xbar_demux;

	component MySoc_rsp_xbar_demux_005 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(92 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component MySoc_rsp_xbar_demux_005;

	component MySoc_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(92 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                        -- ready
			sink4_valid         : in  std_logic                     := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component MySoc_rsp_xbar_mux;

	component MySoc_rsp_xbar_mux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(92 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                        -- ready
			sink4_valid         : in  std_logic                     := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                        -- ready
			sink5_valid         : in  std_logic                     := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                        -- ready
			sink6_valid         : in  std_logic                     := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready         : out std_logic;                                        -- ready
			sink7_valid         : in  std_logic                     := 'X';             -- valid
			sink7_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink7_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink7_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready         : out std_logic;                                        -- ready
			sink8_valid         : in  std_logic                     := 'X';             -- valid
			sink8_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink8_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink8_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready         : out std_logic;                                        -- ready
			sink9_valid         : in  std_logic                     := 'X';             -- valid
			sink9_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink9_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink9_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component MySoc_rsp_xbar_mux_001;

	component MySoc_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component MySoc_irq_mapper;

	component mysoc_nios_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(17 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component mysoc_nios_instruction_master_translator;

	component mysoc_nios_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(17 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component mysoc_nios_data_master_translator;

	component mysoc_nios_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component mysoc_nios_jtag_debug_module_translator;

	component mysoc_ram_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(13 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component mysoc_ram_s1_translator;

	component mysoc_jtag_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component mysoc_jtag_avalon_jtag_slave_translator;

	component mysoc_sysid_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component mysoc_sysid_control_slave_translator;

	component mysoc_performance_counter_0_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(3 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_read                  : out std_logic;                                        -- read
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component mysoc_performance_counter_0_control_slave_translator;

	component mysoc_m_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component mysoc_m_s1_translator;

	component mysoc_res_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component mysoc_res_s1_translator;

	component mysoc_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component mysoc_rst_controller;

	component mysoc_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component mysoc_rst_controller_001;

	signal nios_instruction_master_waitrequest                                                                      : std_logic;                     -- nios_instruction_master_translator:av_waitrequest -> nios:i_waitrequest
	signal nios_instruction_master_address                                                                          : std_logic_vector(17 downto 0); -- nios:i_address -> nios_instruction_master_translator:av_address
	signal nios_instruction_master_read                                                                             : std_logic;                     -- nios:i_read -> nios_instruction_master_translator:av_read
	signal nios_instruction_master_readdata                                                                         : std_logic_vector(31 downto 0); -- nios_instruction_master_translator:av_readdata -> nios:i_readdata
	signal nios_data_master_waitrequest                                                                             : std_logic;                     -- nios_data_master_translator:av_waitrequest -> nios:d_waitrequest
	signal nios_data_master_writedata                                                                               : std_logic_vector(31 downto 0); -- nios:d_writedata -> nios_data_master_translator:av_writedata
	signal nios_data_master_address                                                                                 : std_logic_vector(17 downto 0); -- nios:d_address -> nios_data_master_translator:av_address
	signal nios_data_master_write                                                                                   : std_logic;                     -- nios:d_write -> nios_data_master_translator:av_write
	signal nios_data_master_read                                                                                    : std_logic;                     -- nios:d_read -> nios_data_master_translator:av_read
	signal nios_data_master_readdata                                                                                : std_logic_vector(31 downto 0); -- nios_data_master_translator:av_readdata -> nios:d_readdata
	signal nios_data_master_debugaccess                                                                             : std_logic;                     -- nios:jtag_debug_module_debugaccess_to_roms -> nios_data_master_translator:av_debugaccess
	signal nios_data_master_byteenable                                                                              : std_logic_vector(3 downto 0);  -- nios:d_byteenable -> nios_data_master_translator:av_byteenable
	signal nios_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                                        : std_logic;                     -- nios:jtag_debug_module_waitrequest -> nios_jtag_debug_module_translator:av_waitrequest
	signal nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                          : std_logic_vector(31 downto 0); -- nios_jtag_debug_module_translator:av_writedata -> nios:jtag_debug_module_writedata
	signal nios_jtag_debug_module_translator_avalon_anti_slave_0_address                                            : std_logic_vector(8 downto 0);  -- nios_jtag_debug_module_translator:av_address -> nios:jtag_debug_module_address
	signal nios_jtag_debug_module_translator_avalon_anti_slave_0_write                                              : std_logic;                     -- nios_jtag_debug_module_translator:av_write -> nios:jtag_debug_module_write
	signal nios_jtag_debug_module_translator_avalon_anti_slave_0_read                                               : std_logic;                     -- nios_jtag_debug_module_translator:av_read -> nios:jtag_debug_module_read
	signal nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                           : std_logic_vector(31 downto 0); -- nios:jtag_debug_module_readdata -> nios_jtag_debug_module_translator:av_readdata
	signal nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                        : std_logic;                     -- nios_jtag_debug_module_translator:av_debugaccess -> nios:jtag_debug_module_debugaccess
	signal nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                         : std_logic_vector(3 downto 0);  -- nios_jtag_debug_module_translator:av_byteenable -> nios:jtag_debug_module_byteenable
	signal ram_s1_translator_avalon_anti_slave_0_writedata                                                          : std_logic_vector(31 downto 0); -- ram_s1_translator:av_writedata -> ram:writedata
	signal ram_s1_translator_avalon_anti_slave_0_address                                                            : std_logic_vector(13 downto 0); -- ram_s1_translator:av_address -> ram:address
	signal ram_s1_translator_avalon_anti_slave_0_chipselect                                                         : std_logic;                     -- ram_s1_translator:av_chipselect -> ram:chipselect
	signal ram_s1_translator_avalon_anti_slave_0_clken                                                              : std_logic;                     -- ram_s1_translator:av_clken -> ram:clken
	signal ram_s1_translator_avalon_anti_slave_0_write                                                              : std_logic;                     -- ram_s1_translator:av_write -> ram:write
	signal ram_s1_translator_avalon_anti_slave_0_readdata                                                           : std_logic_vector(31 downto 0); -- ram:readdata -> ram_s1_translator:av_readdata
	signal ram_s1_translator_avalon_anti_slave_0_byteenable                                                         : std_logic_vector(3 downto 0);  -- ram_s1_translator:av_byteenable -> ram:byteenable
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                                        : std_logic;                     -- jtag:av_waitrequest -> jtag_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                          : std_logic_vector(31 downto 0); -- jtag_avalon_jtag_slave_translator:av_writedata -> jtag:av_writedata
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                            : std_logic_vector(0 downto 0);  -- jtag_avalon_jtag_slave_translator:av_address -> jtag:av_address
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                                         : std_logic;                     -- jtag_avalon_jtag_slave_translator:av_chipselect -> jtag:av_chipselect
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                              : std_logic;                     -- jtag_avalon_jtag_slave_translator:av_write -> jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                               : std_logic;                     -- jtag_avalon_jtag_slave_translator:av_read -> jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                           : std_logic_vector(31 downto 0); -- jtag:av_readdata -> jtag_avalon_jtag_slave_translator:av_readdata
	signal sysid_control_slave_translator_avalon_anti_slave_0_address                                               : std_logic_vector(0 downto 0);  -- sysid_control_slave_translator:av_address -> sysid:address
	signal sysid_control_slave_translator_avalon_anti_slave_0_readdata                                              : std_logic_vector(31 downto 0); -- sysid:readdata -> sysid_control_slave_translator:av_readdata
	signal performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- performance_counter_0_control_slave_translator:av_writedata -> performance_counter_0:writedata
	signal performance_counter_0_control_slave_translator_avalon_anti_slave_0_address                               : std_logic_vector(3 downto 0);  -- performance_counter_0_control_slave_translator:av_address -> performance_counter_0:address
	signal performance_counter_0_control_slave_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- performance_counter_0_control_slave_translator:av_write -> performance_counter_0:write
	signal performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- performance_counter_0:readdata -> performance_counter_0_control_slave_translator:av_readdata
	signal performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer                         : std_logic;                     -- performance_counter_0_control_slave_translator:av_begintransfer -> performance_counter_0:begintransfer
	signal m_s1_translator_avalon_anti_slave_0_writedata                                                            : std_logic_vector(31 downto 0); -- m_s1_translator:av_writedata -> m:writedata
	signal m_s1_translator_avalon_anti_slave_0_address                                                              : std_logic_vector(1 downto 0);  -- m_s1_translator:av_address -> m:address
	signal m_s1_translator_avalon_anti_slave_0_chipselect                                                           : std_logic;                     -- m_s1_translator:av_chipselect -> m:chipselect
	signal m_s1_translator_avalon_anti_slave_0_write                                                                : std_logic;                     -- m_s1_translator:av_write -> m_s1_translator_avalon_anti_slave_0_write:in
	signal m_s1_translator_avalon_anti_slave_0_readdata                                                             : std_logic_vector(31 downto 0); -- m:readdata -> m_s1_translator:av_readdata
	signal mult_s1_translator_avalon_anti_slave_0_writedata                                                         : std_logic_vector(31 downto 0); -- mult_s1_translator:av_writedata -> mult:writedata
	signal mult_s1_translator_avalon_anti_slave_0_address                                                           : std_logic_vector(1 downto 0);  -- mult_s1_translator:av_address -> mult:address
	signal mult_s1_translator_avalon_anti_slave_0_chipselect                                                        : std_logic;                     -- mult_s1_translator:av_chipselect -> mult:chipselect
	signal mult_s1_translator_avalon_anti_slave_0_write                                                             : std_logic;                     -- mult_s1_translator:av_write -> mult_s1_translator_avalon_anti_slave_0_write:in
	signal mult_s1_translator_avalon_anti_slave_0_readdata                                                          : std_logic_vector(31 downto 0); -- mult:readdata -> mult_s1_translator:av_readdata
	signal res_s1_translator_avalon_anti_slave_0_address                                                            : std_logic_vector(1 downto 0);  -- res_s1_translator:av_address -> res:address
	signal res_s1_translator_avalon_anti_slave_0_readdata                                                           : std_logic_vector(31 downto 0); -- res:readdata -> res_s1_translator:av_readdata
	signal prt_s1_translator_avalon_anti_slave_0_address                                                            : std_logic_vector(1 downto 0);  -- prt_s1_translator:av_address -> prt:address
	signal prt_s1_translator_avalon_anti_slave_0_readdata                                                           : std_logic_vector(31 downto 0); -- prt:readdata -> prt_s1_translator:av_readdata
	signal go_s1_translator_avalon_anti_slave_0_writedata                                                           : std_logic_vector(31 downto 0); -- go_s1_translator:av_writedata -> go:writedata
	signal go_s1_translator_avalon_anti_slave_0_address                                                             : std_logic_vector(1 downto 0);  -- go_s1_translator:av_address -> go:address
	signal go_s1_translator_avalon_anti_slave_0_chipselect                                                          : std_logic;                     -- go_s1_translator:av_chipselect -> go:chipselect
	signal go_s1_translator_avalon_anti_slave_0_write                                                               : std_logic;                     -- go_s1_translator:av_write -> go_s1_translator_avalon_anti_slave_0_write:in
	signal go_s1_translator_avalon_anti_slave_0_readdata                                                            : std_logic_vector(31 downto 0); -- go:readdata -> go_s1_translator:av_readdata
	signal nios_instruction_master_translator_avalon_universal_master_0_waitrequest                                 : std_logic;                     -- nios_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios_instruction_master_translator:uav_waitrequest
	signal nios_instruction_master_translator_avalon_universal_master_0_burstcount                                  : std_logic_vector(2 downto 0);  -- nios_instruction_master_translator:uav_burstcount -> nios_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios_instruction_master_translator_avalon_universal_master_0_writedata                                   : std_logic_vector(31 downto 0); -- nios_instruction_master_translator:uav_writedata -> nios_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios_instruction_master_translator_avalon_universal_master_0_address                                     : std_logic_vector(17 downto 0); -- nios_instruction_master_translator:uav_address -> nios_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios_instruction_master_translator_avalon_universal_master_0_lock                                        : std_logic;                     -- nios_instruction_master_translator:uav_lock -> nios_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios_instruction_master_translator_avalon_universal_master_0_write                                       : std_logic;                     -- nios_instruction_master_translator:uav_write -> nios_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios_instruction_master_translator_avalon_universal_master_0_read                                        : std_logic;                     -- nios_instruction_master_translator:uav_read -> nios_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios_instruction_master_translator_avalon_universal_master_0_readdata                                    : std_logic_vector(31 downto 0); -- nios_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios_instruction_master_translator:uav_readdata
	signal nios_instruction_master_translator_avalon_universal_master_0_debugaccess                                 : std_logic;                     -- nios_instruction_master_translator:uav_debugaccess -> nios_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios_instruction_master_translator_avalon_universal_master_0_byteenable                                  : std_logic_vector(3 downto 0);  -- nios_instruction_master_translator:uav_byteenable -> nios_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios_instruction_master_translator_avalon_universal_master_0_readdatavalid                               : std_logic;                     -- nios_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios_instruction_master_translator:uav_readdatavalid
	signal nios_data_master_translator_avalon_universal_master_0_waitrequest                                        : std_logic;                     -- nios_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios_data_master_translator:uav_waitrequest
	signal nios_data_master_translator_avalon_universal_master_0_burstcount                                         : std_logic_vector(2 downto 0);  -- nios_data_master_translator:uav_burstcount -> nios_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios_data_master_translator_avalon_universal_master_0_writedata                                          : std_logic_vector(31 downto 0); -- nios_data_master_translator:uav_writedata -> nios_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios_data_master_translator_avalon_universal_master_0_address                                            : std_logic_vector(17 downto 0); -- nios_data_master_translator:uav_address -> nios_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios_data_master_translator_avalon_universal_master_0_lock                                               : std_logic;                     -- nios_data_master_translator:uav_lock -> nios_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios_data_master_translator_avalon_universal_master_0_write                                              : std_logic;                     -- nios_data_master_translator:uav_write -> nios_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios_data_master_translator_avalon_universal_master_0_read                                               : std_logic;                     -- nios_data_master_translator:uav_read -> nios_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios_data_master_translator_avalon_universal_master_0_readdata                                           : std_logic_vector(31 downto 0); -- nios_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios_data_master_translator:uav_readdata
	signal nios_data_master_translator_avalon_universal_master_0_debugaccess                                        : std_logic;                     -- nios_data_master_translator:uav_debugaccess -> nios_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios_data_master_translator_avalon_universal_master_0_byteenable                                         : std_logic_vector(3 downto 0);  -- nios_data_master_translator:uav_byteenable -> nios_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios_data_master_translator_avalon_universal_master_0_readdatavalid                                      : std_logic;                     -- nios_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios_data_master_translator:uav_readdatavalid
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                          : std_logic;                     -- nios_jtag_debug_module_translator:uav_waitrequest -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                           : std_logic_vector(2 downto 0);  -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios_jtag_debug_module_translator:uav_burstcount
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                            : std_logic_vector(31 downto 0); -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios_jtag_debug_module_translator:uav_writedata
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                              : std_logic_vector(17 downto 0); -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios_jtag_debug_module_translator:uav_address
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                                : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios_jtag_debug_module_translator:uav_write
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                                 : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios_jtag_debug_module_translator:uav_lock
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                                 : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios_jtag_debug_module_translator:uav_read
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                             : std_logic_vector(31 downto 0); -- nios_jtag_debug_module_translator:uav_readdata -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                        : std_logic;                     -- nios_jtag_debug_module_translator:uav_readdatavalid -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                          : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios_jtag_debug_module_translator:uav_debugaccess
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                           : std_logic_vector(3 downto 0);  -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios_jtag_debug_module_translator:uav_byteenable
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                   : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                         : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                 : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                          : std_logic_vector(93 downto 0); -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                         : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                      : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket              : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                       : std_logic_vector(93 downto 0); -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                      : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                    : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                     : std_logic_vector(33 downto 0); -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                    : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                          : std_logic;                     -- ram_s1_translator:uav_waitrequest -> ram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                           : std_logic_vector(2 downto 0);  -- ram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ram_s1_translator:uav_burstcount
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                            : std_logic_vector(31 downto 0); -- ram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ram_s1_translator:uav_writedata
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_address                                              : std_logic_vector(17 downto 0); -- ram_s1_translator_avalon_universal_slave_0_agent:m0_address -> ram_s1_translator:uav_address
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_write                                                : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:m0_write -> ram_s1_translator:uav_write
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                 : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ram_s1_translator:uav_lock
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_read                                                 : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:m0_read -> ram_s1_translator:uav_read
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                             : std_logic_vector(31 downto 0); -- ram_s1_translator:uav_readdata -> ram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                        : std_logic;                     -- ram_s1_translator:uav_readdatavalid -> ram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                          : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ram_s1_translator:uav_debugaccess
	signal ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                           : std_logic_vector(3 downto 0);  -- ram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ram_s1_translator:uav_byteenable
	signal ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                   : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                         : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                 : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                          : std_logic_vector(93 downto 0); -- ram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                         : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                      : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                              : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                       : std_logic_vector(93 downto 0); -- ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                      : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                    : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                     : std_logic_vector(33 downto 0); -- ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                    : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                          : std_logic;                     -- jtag_avalon_jtag_slave_translator:uav_waitrequest -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                           : std_logic_vector(2 downto 0);  -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                            : std_logic_vector(31 downto 0); -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_avalon_jtag_slave_translator:uav_writedata
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                              : std_logic_vector(17 downto 0); -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_avalon_jtag_slave_translator:uav_address
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                                : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_avalon_jtag_slave_translator:uav_write
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                                 : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_avalon_jtag_slave_translator:uav_lock
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                                 : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_avalon_jtag_slave_translator:uav_read
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                             : std_logic_vector(31 downto 0); -- jtag_avalon_jtag_slave_translator:uav_readdata -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                        : std_logic;                     -- jtag_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                          : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                           : std_logic_vector(3 downto 0);  -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                   : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                         : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                 : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                          : std_logic_vector(93 downto 0); -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                         : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                      : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket              : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                       : std_logic_vector(93 downto 0); -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                      : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                    : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                     : std_logic_vector(33 downto 0); -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                    : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                             : std_logic;                     -- sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                              : std_logic_vector(2 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                               : std_logic_vector(31 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                 : std_logic_vector(17 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                   : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                    : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                    : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                : std_logic_vector(31 downto 0); -- sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                           : std_logic;                     -- sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                             : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                              : std_logic_vector(3 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                      : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                            : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                    : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                             : std_logic_vector(93 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                            : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                   : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                         : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                 : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                          : std_logic_vector(93 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                         : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                       : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                        : std_logic_vector(33 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                       : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- performance_counter_0_control_slave_translator:uav_waitrequest -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_0_control_slave_translator:uav_burstcount
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_0_control_slave_translator:uav_writedata
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(17 downto 0); -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_0_control_slave_translator:uav_address
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_0_control_slave_translator:uav_write
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_0_control_slave_translator:uav_lock
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_0_control_slave_translator:uav_read
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- performance_counter_0_control_slave_translator:uav_readdata -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- performance_counter_0_control_slave_translator:uav_readdatavalid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_0_control_slave_translator:uav_debugaccess
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_0_control_slave_translator:uav_byteenable
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(93 downto 0); -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(93 downto 0); -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0); -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                            : std_logic;                     -- m_s1_translator:uav_waitrequest -> m_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                             : std_logic_vector(2 downto 0);  -- m_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> m_s1_translator:uav_burstcount
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                              : std_logic_vector(31 downto 0); -- m_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> m_s1_translator:uav_writedata
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_address                                                : std_logic_vector(17 downto 0); -- m_s1_translator_avalon_universal_slave_0_agent:m0_address -> m_s1_translator:uav_address
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_write                                                  : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:m0_write -> m_s1_translator:uav_write
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                   : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:m0_lock -> m_s1_translator:uav_lock
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_read                                                   : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:m0_read -> m_s1_translator:uav_read
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                               : std_logic_vector(31 downto 0); -- m_s1_translator:uav_readdata -> m_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                          : std_logic;                     -- m_s1_translator:uav_readdatavalid -> m_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                            : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> m_s1_translator:uav_debugaccess
	signal m_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                             : std_logic_vector(3 downto 0);  -- m_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> m_s1_translator:uav_byteenable
	signal m_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                     : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal m_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                           : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal m_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                   : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal m_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                            : std_logic_vector(93 downto 0); -- m_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal m_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                           : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> m_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                  : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> m_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                        : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> m_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                                : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> m_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                         : std_logic_vector(93 downto 0); -- m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> m_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                        : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                      : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> m_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                       : std_logic_vector(33 downto 0); -- m_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> m_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                      : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> m_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                         : std_logic;                     -- mult_s1_translator:uav_waitrequest -> mult_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                          : std_logic_vector(2 downto 0);  -- mult_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mult_s1_translator:uav_burstcount
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                           : std_logic_vector(31 downto 0); -- mult_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mult_s1_translator:uav_writedata
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_address                                             : std_logic_vector(17 downto 0); -- mult_s1_translator_avalon_universal_slave_0_agent:m0_address -> mult_s1_translator:uav_address
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_write                                               : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:m0_write -> mult_s1_translator:uav_write
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mult_s1_translator:uav_lock
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_read                                                : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:m0_read -> mult_s1_translator:uav_read
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                            : std_logic_vector(31 downto 0); -- mult_s1_translator:uav_readdata -> mult_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                       : std_logic;                     -- mult_s1_translator:uav_readdatavalid -> mult_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                         : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mult_s1_translator:uav_debugaccess
	signal mult_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                          : std_logic_vector(3 downto 0);  -- mult_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mult_s1_translator:uav_byteenable
	signal mult_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                  : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal mult_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                        : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal mult_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal mult_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                         : std_logic_vector(93 downto 0); -- mult_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal mult_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                        : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mult_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                               : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mult_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                     : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mult_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                             : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mult_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                      : std_logic_vector(93 downto 0); -- mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mult_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                     : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                   : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mult_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                    : std_logic_vector(33 downto 0); -- mult_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mult_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                   : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mult_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                          : std_logic;                     -- res_s1_translator:uav_waitrequest -> res_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                           : std_logic_vector(2 downto 0);  -- res_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> res_s1_translator:uav_burstcount
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                            : std_logic_vector(31 downto 0); -- res_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> res_s1_translator:uav_writedata
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_address                                              : std_logic_vector(17 downto 0); -- res_s1_translator_avalon_universal_slave_0_agent:m0_address -> res_s1_translator:uav_address
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_write                                                : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:m0_write -> res_s1_translator:uav_write
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                 : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:m0_lock -> res_s1_translator:uav_lock
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_read                                                 : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:m0_read -> res_s1_translator:uav_read
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                             : std_logic_vector(31 downto 0); -- res_s1_translator:uav_readdata -> res_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                        : std_logic;                     -- res_s1_translator:uav_readdatavalid -> res_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                          : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> res_s1_translator:uav_debugaccess
	signal res_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                           : std_logic_vector(3 downto 0);  -- res_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> res_s1_translator:uav_byteenable
	signal res_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                   : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal res_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                         : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal res_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                 : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal res_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                          : std_logic_vector(93 downto 0); -- res_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal res_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                         : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> res_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> res_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                      : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> res_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                              : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> res_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                       : std_logic_vector(93 downto 0); -- res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> res_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                      : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                    : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> res_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                     : std_logic_vector(33 downto 0); -- res_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> res_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                    : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> res_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                          : std_logic;                     -- prt_s1_translator:uav_waitrequest -> prt_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                           : std_logic_vector(2 downto 0);  -- prt_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> prt_s1_translator:uav_burstcount
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                            : std_logic_vector(31 downto 0); -- prt_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> prt_s1_translator:uav_writedata
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_address                                              : std_logic_vector(17 downto 0); -- prt_s1_translator_avalon_universal_slave_0_agent:m0_address -> prt_s1_translator:uav_address
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_write                                                : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:m0_write -> prt_s1_translator:uav_write
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                 : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:m0_lock -> prt_s1_translator:uav_lock
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_read                                                 : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:m0_read -> prt_s1_translator:uav_read
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                             : std_logic_vector(31 downto 0); -- prt_s1_translator:uav_readdata -> prt_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                        : std_logic;                     -- prt_s1_translator:uav_readdatavalid -> prt_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                          : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> prt_s1_translator:uav_debugaccess
	signal prt_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                           : std_logic_vector(3 downto 0);  -- prt_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> prt_s1_translator:uav_byteenable
	signal prt_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                   : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal prt_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                         : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal prt_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                 : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal prt_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                          : std_logic_vector(93 downto 0); -- prt_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal prt_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                         : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> prt_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> prt_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                      : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> prt_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                              : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> prt_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                       : std_logic_vector(93 downto 0); -- prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> prt_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                      : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                    : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> prt_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                     : std_logic_vector(33 downto 0); -- prt_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> prt_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                    : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> prt_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                           : std_logic;                     -- go_s1_translator:uav_waitrequest -> go_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                            : std_logic_vector(2 downto 0);  -- go_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> go_s1_translator:uav_burstcount
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                             : std_logic_vector(31 downto 0); -- go_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> go_s1_translator:uav_writedata
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_address                                               : std_logic_vector(17 downto 0); -- go_s1_translator_avalon_universal_slave_0_agent:m0_address -> go_s1_translator:uav_address
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_write                                                 : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:m0_write -> go_s1_translator:uav_write
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                  : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:m0_lock -> go_s1_translator:uav_lock
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_read                                                  : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:m0_read -> go_s1_translator:uav_read
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                              : std_logic_vector(31 downto 0); -- go_s1_translator:uav_readdata -> go_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                         : std_logic;                     -- go_s1_translator:uav_readdatavalid -> go_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                           : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> go_s1_translator:uav_debugaccess
	signal go_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                            : std_logic_vector(3 downto 0);  -- go_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> go_s1_translator:uav_byteenable
	signal go_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                    : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal go_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                          : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal go_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                  : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal go_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                           : std_logic_vector(93 downto 0); -- go_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal go_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                          : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> go_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                 : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> go_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                       : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> go_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                               : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> go_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                        : std_logic_vector(93 downto 0); -- go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> go_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                       : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                     : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> go_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                      : std_logic_vector(33 downto 0); -- go_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> go_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                     : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> go_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                        : std_logic;                     -- nios_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                              : std_logic;                     -- nios_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket                      : std_logic;                     -- nios_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data                               : std_logic_vector(92 downto 0); -- nios_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                              : std_logic;                     -- addr_router:sink_ready -> nios_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                               : std_logic;                     -- nios_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios_data_master_translator_avalon_universal_master_0_agent_cp_valid                                     : std_logic;                     -- nios_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                             : std_logic;                     -- nios_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios_data_master_translator_avalon_universal_master_0_agent_cp_data                                      : std_logic_vector(92 downto 0); -- nios_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios_data_master_translator_avalon_universal_master_0_agent_cp_ready                                     : std_logic;                     -- addr_router_001:sink_ready -> nios_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                          : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                                : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                        : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                                 : std_logic_vector(92 downto 0); -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                                : std_logic;                     -- id_router:sink_ready -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                          : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal ram_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                        : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal ram_s1_translator_avalon_universal_slave_0_agent_rp_data                                                 : std_logic_vector(92 downto 0); -- ram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal ram_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                : std_logic;                     -- id_router_001:sink_ready -> ram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                          : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                                : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                        : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                                 : std_logic_vector(92 downto 0); -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                                : std_logic;                     -- id_router_002:sink_ready -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                             : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                   : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                           : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                    : std_logic_vector(92 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                   : std_logic;                     -- id_router_003:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(92 downto 0); -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router_004:sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal m_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                            : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal m_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                  : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal m_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                          : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal m_s1_translator_avalon_universal_slave_0_agent_rp_data                                                   : std_logic_vector(92 downto 0); -- m_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal m_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                  : std_logic;                     -- id_router_005:sink_ready -> m_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal mult_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                         : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal mult_s1_translator_avalon_universal_slave_0_agent_rp_valid                                               : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal mult_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                       : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal mult_s1_translator_avalon_universal_slave_0_agent_rp_data                                                : std_logic_vector(92 downto 0); -- mult_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal mult_s1_translator_avalon_universal_slave_0_agent_rp_ready                                               : std_logic;                     -- id_router_006:sink_ready -> mult_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal res_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                          : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal res_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal res_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                        : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal res_s1_translator_avalon_universal_slave_0_agent_rp_data                                                 : std_logic_vector(92 downto 0); -- res_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal res_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                : std_logic;                     -- id_router_007:sink_ready -> res_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal prt_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                          : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal prt_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal prt_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                        : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal prt_s1_translator_avalon_universal_slave_0_agent_rp_data                                                 : std_logic_vector(92 downto 0); -- prt_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal prt_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                : std_logic;                     -- id_router_008:sink_ready -> prt_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal go_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                           : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal go_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                 : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal go_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                         : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal go_s1_translator_avalon_universal_slave_0_agent_rp_data                                                  : std_logic_vector(92 downto 0); -- go_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal go_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                 : std_logic;                     -- id_router_009:sink_ready -> go_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal rst_controller_reset_out_reset                                                                           : std_logic;                     -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, id_router:reset, irq_mapper:reset, nios_data_master_translator:reset, nios_data_master_translator_avalon_universal_master_0_agent:reset, nios_instruction_master_translator:reset, nios_instruction_master_translator_avalon_universal_master_0_agent:reset, nios_jtag_debug_module_translator:reset, nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                                                                       : std_logic;                     -- rst_controller_001:reset_out -> [cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, go_s1_translator:reset, go_s1_translator_avalon_universal_slave_0_agent:reset, go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, jtag_avalon_jtag_slave_translator:reset, jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, m_s1_translator:reset, m_s1_translator_avalon_universal_slave_0_agent:reset, m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mult_s1_translator:reset, mult_s1_translator_avalon_universal_slave_0_agent:reset, mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, performance_counter_0_control_slave_translator:reset, performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, prt_s1_translator:reset, prt_s1_translator_avalon_universal_slave_0_agent:reset, prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ram:reset, ram_s1_translator:reset, ram_s1_translator_avalon_universal_slave_0_agent:reset, ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, res_s1_translator:reset, res_s1_translator_avalon_universal_slave_0_agent:reset, res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rst_controller_001_reset_out_reset:in, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal rst_controller_001_reset_out_reset_req                                                                   : std_logic;                     -- rst_controller_001:reset_req -> ram:reset_req
	signal nios_jtag_debug_module_reset_reset                                                                       : std_logic;                     -- nios:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1
	signal cmd_xbar_demux_src0_endofpacket                                                                          : std_logic;                     -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                                : std_logic;                     -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                                 : std_logic_vector(92 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                              : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                                : std_logic;                     -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                          : std_logic;                     -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                                : std_logic;                     -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                                 : std_logic_vector(92 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                              : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                                : std_logic;                     -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                          : std_logic;                     -- cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                                : std_logic;                     -- cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal cmd_xbar_demux_src2_data                                                                                 : std_logic_vector(92 downto 0); -- cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	signal cmd_xbar_demux_src2_channel                                                                              : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_src2_ready                                                                                : std_logic;                     -- cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	signal cmd_xbar_demux_src3_endofpacket                                                                          : std_logic;                     -- cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                                : std_logic;                     -- cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal cmd_xbar_demux_src3_data                                                                                 : std_logic_vector(92 downto 0); -- cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	signal cmd_xbar_demux_src3_channel                                                                              : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_src3_ready                                                                                : std_logic;                     -- cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	signal cmd_xbar_demux_src4_endofpacket                                                                          : std_logic;                     -- cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	signal cmd_xbar_demux_src4_valid                                                                                : std_logic;                     -- cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	signal cmd_xbar_demux_src4_startofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	signal cmd_xbar_demux_src4_data                                                                                 : std_logic_vector(92 downto 0); -- cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	signal cmd_xbar_demux_src4_channel                                                                              : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	signal cmd_xbar_demux_src4_ready                                                                                : std_logic;                     -- cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                            : std_logic;                     -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                            : std_logic;                     -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                            : std_logic;                     -- cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal cmd_xbar_demux_001_src3_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	signal cmd_xbar_demux_001_src3_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_001_src3_ready                                                                            : std_logic;                     -- cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	signal cmd_xbar_demux_001_src4_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	signal cmd_xbar_demux_001_src4_ready                                                                            : std_logic;                     -- cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	signal cmd_xbar_demux_001_src5_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src5_endofpacket -> m_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src5_valid -> m_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src5_startofpacket -> m_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src5_data -> m_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src5_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src5_channel -> m_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src6_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src6_endofpacket -> mult_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src6_valid -> mult_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src6_startofpacket -> mult_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src6_data -> mult_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src6_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src6_channel -> mult_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src7_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src7_endofpacket -> res_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src7_valid -> res_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src7_startofpacket -> res_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src7_data -> res_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src7_channel -> res_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src8_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src8_endofpacket -> prt_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src8_valid -> prt_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src8_startofpacket -> prt_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src8_data -> prt_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src8_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src8_channel -> prt_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src9_endofpacket                                                                      : std_logic;                     -- cmd_xbar_demux_001:src9_endofpacket -> go_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                            : std_logic;                     -- cmd_xbar_demux_001:src9_valid -> go_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                                    : std_logic;                     -- cmd_xbar_demux_001:src9_startofpacket -> go_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                             : std_logic_vector(92 downto 0); -- cmd_xbar_demux_001:src9_data -> go_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src9_channel                                                                          : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src9_channel -> go_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                          : std_logic;                     -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                                : std_logic;                     -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                        : std_logic;                     -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                                 : std_logic_vector(92 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                              : std_logic_vector(9 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                                : std_logic;                     -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                          : std_logic;                     -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                                : std_logic;                     -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                        : std_logic;                     -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                                 : std_logic_vector(92 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                              : std_logic_vector(9 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                                : std_logic;                     -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                            : std_logic;                     -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_002_src1_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                            : std_logic;                     -- rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src1_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src1_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_003_src1_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                            : std_logic;                     -- rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src1_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src1_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_004_src1_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src1_valid                                                                            : std_logic;                     -- rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src1_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src1_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src1_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src1_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                      : std_logic;                     -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                            : std_logic;                     -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                             : std_logic_vector(92 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                          : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                            : std_logic;                     -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal addr_router_src_endofpacket                                                                              : std_logic;                     -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                                    : std_logic;                     -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                            : std_logic;                     -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                     : std_logic_vector(92 downto 0); -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                                  : std_logic_vector(9 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                                    : std_logic;                     -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                             : std_logic;                     -- rsp_xbar_mux:src_endofpacket -> nios_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                   : std_logic;                     -- rsp_xbar_mux:src_valid -> nios_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                           : std_logic;                     -- rsp_xbar_mux:src_startofpacket -> nios_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                                    : std_logic_vector(92 downto 0); -- rsp_xbar_mux:src_data -> nios_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                                 : std_logic_vector(9 downto 0);  -- rsp_xbar_mux:src_channel -> nios_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                                   : std_logic;                     -- nios_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                          : std_logic;                     -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                                : std_logic;                     -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                        : std_logic;                     -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                                 : std_logic_vector(92 downto 0); -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                              : std_logic_vector(9 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                                : std_logic;                     -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                         : std_logic;                     -- rsp_xbar_mux_001:src_endofpacket -> nios_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                               : std_logic;                     -- rsp_xbar_mux_001:src_valid -> nios_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                       : std_logic;                     -- rsp_xbar_mux_001:src_startofpacket -> nios_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                                : std_logic_vector(92 downto 0); -- rsp_xbar_mux_001:src_data -> nios_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                             : std_logic_vector(9 downto 0);  -- rsp_xbar_mux_001:src_channel -> nios_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                               : std_logic;                     -- nios_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                             : std_logic;                     -- cmd_xbar_mux:src_endofpacket -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                   : std_logic;                     -- cmd_xbar_mux:src_valid -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                           : std_logic;                     -- cmd_xbar_mux:src_startofpacket -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                    : std_logic_vector(92 downto 0); -- cmd_xbar_mux:src_data -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                                 : std_logic_vector(9 downto 0);  -- cmd_xbar_mux:src_channel -> nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                   : std_logic;                     -- nios_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                                : std_logic;                     -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                      : std_logic;                     -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                              : std_logic;                     -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                       : std_logic_vector(92 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                    : std_logic_vector(9 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                      : std_logic;                     -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                         : std_logic;                     -- cmd_xbar_mux_001:src_endofpacket -> ram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                               : std_logic;                     -- cmd_xbar_mux_001:src_valid -> ram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                       : std_logic;                     -- cmd_xbar_mux_001:src_startofpacket -> ram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                                : std_logic_vector(92 downto 0); -- cmd_xbar_mux_001:src_data -> ram_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                             : std_logic_vector(9 downto 0);  -- cmd_xbar_mux_001:src_channel -> ram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                               : std_logic;                     -- ram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                            : std_logic;                     -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                                  : std_logic;                     -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                          : std_logic;                     -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                                         : std_logic;                     -- cmd_xbar_mux_002:src_endofpacket -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                               : std_logic;                     -- cmd_xbar_mux_002:src_valid -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                                       : std_logic;                     -- cmd_xbar_mux_002:src_startofpacket -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                                : std_logic_vector(92 downto 0); -- cmd_xbar_mux_002:src_data -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_002_src_channel                                                                             : std_logic_vector(9 downto 0);  -- cmd_xbar_mux_002:src_channel -> jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_002_src_ready                                                                               : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	signal id_router_002_src_endofpacket                                                                            : std_logic;                     -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                                  : std_logic;                     -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                          : std_logic;                     -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_mux_003_src_endofpacket                                                                         : std_logic;                     -- cmd_xbar_mux_003:src_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                               : std_logic;                     -- cmd_xbar_mux_003:src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                       : std_logic;                     -- cmd_xbar_mux_003:src_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                                : std_logic_vector(92 downto 0); -- cmd_xbar_mux_003:src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_003_src_channel                                                                             : std_logic_vector(9 downto 0);  -- cmd_xbar_mux_003:src_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_003_src_ready                                                                               : std_logic;                     -- sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	signal id_router_003_src_endofpacket                                                                            : std_logic;                     -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                                  : std_logic;                     -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                          : std_logic;                     -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_mux_004_src_endofpacket                                                                         : std_logic;                     -- cmd_xbar_mux_004:src_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_004_src_valid                                                                               : std_logic;                     -- cmd_xbar_mux_004:src_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_004_src_startofpacket                                                                       : std_logic;                     -- cmd_xbar_mux_004:src_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_004_src_data                                                                                : std_logic_vector(92 downto 0); -- cmd_xbar_mux_004:src_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_004_src_channel                                                                             : std_logic_vector(9 downto 0);  -- cmd_xbar_mux_004:src_channel -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_004_src_ready                                                                               : std_logic;                     -- performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	signal id_router_004_src_endofpacket                                                                            : std_logic;                     -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                                  : std_logic;                     -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                          : std_logic;                     -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_001_src5_ready                                                                            : std_logic;                     -- m_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	signal id_router_005_src_endofpacket                                                                            : std_logic;                     -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                                  : std_logic;                     -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                          : std_logic;                     -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_001_src6_ready                                                                            : std_logic;                     -- mult_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	signal id_router_006_src_endofpacket                                                                            : std_logic;                     -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                                  : std_logic;                     -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                          : std_logic;                     -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                            : std_logic;                     -- res_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                            : std_logic;                     -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                                  : std_logic;                     -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                          : std_logic;                     -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_001_src8_ready                                                                            : std_logic;                     -- prt_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	signal id_router_008_src_endofpacket                                                                            : std_logic;                     -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                                  : std_logic;                     -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                          : std_logic;                     -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_001_src9_ready                                                                            : std_logic;                     -- go_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	signal id_router_009_src_endofpacket                                                                            : std_logic;                     -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                                  : std_logic;                     -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                          : std_logic;                     -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                                   : std_logic_vector(92 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                                : std_logic_vector(9 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                                  : std_logic;                     -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal irq_mapper_receiver0_irq                                                                                 : std_logic;                     -- jtag:av_irq -> irq_mapper:receiver0_irq
	signal nios_d_irq_irq                                                                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios:d_irq
	signal reset_reset_n_ports_inv                                                                                  : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                                    : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag:av_write_n
	signal jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                                     : std_logic;                     -- jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag:av_read_n
	signal m_s1_translator_avalon_anti_slave_0_write_ports_inv                                                      : std_logic;                     -- m_s1_translator_avalon_anti_slave_0_write:inv -> m:write_n
	signal mult_s1_translator_avalon_anti_slave_0_write_ports_inv                                                   : std_logic;                     -- mult_s1_translator_avalon_anti_slave_0_write:inv -> mult:write_n
	signal go_s1_translator_avalon_anti_slave_0_write_ports_inv                                                     : std_logic;                     -- go_s1_translator_avalon_anti_slave_0_write:inv -> go:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> nios:reset_n
	signal rst_controller_001_reset_out_reset_ports_inv                                                             : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [go:reset_n, jtag:rst_n, m:reset_n, mult:reset_n, performance_counter_0:reset_n, prt:reset_n, res:reset_n, sysid:reset_n]

begin

	nios : component MySoc_nios
		port map (
			clk                                   => clk_clk,                                                           --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                          --                   reset_n.reset_n
			d_address                             => nios_data_master_address,                                          --               data_master.address
			d_byteenable                          => nios_data_master_byteenable,                                       --                          .byteenable
			d_read                                => nios_data_master_read,                                             --                          .read
			d_readdata                            => nios_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => nios_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => nios_data_master_write,                                            --                          .write
			d_writedata                           => nios_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => nios_instruction_master_address,                                   --        instruction_master.address
			i_read                                => nios_instruction_master_read,                                      --                          .read
			i_readdata                            => nios_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => nios_instruction_master_waitrequest,                               --                          .waitrequest
			d_irq                                 => nios_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios_jtag_debug_module_reset_reset,                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => nios_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => nios_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => nios_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                               -- custom_instruction_master.readra
		);

	ram : component MySoc_ram
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => ram_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => ram_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => ram_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => ram_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => ram_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => ram_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => ram_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req            --       .reset_req
		);

	jtag : component MySoc_jtag
		port map (
			clk            => clk_clk,                                                               --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                          --             reset.reset_n
			av_chipselect  => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                               --               irq.irq
		);

	sysid : component MySoc_sysid
		port map (
			clock    => clk_clk,                                                       --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,                  --         reset.reset_n
			readdata => sysid_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	m : component MySoc_m
		port map (
			clk        => clk_clk,                                             --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => m_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => m_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => m_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => m_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => m_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => m_export                                             -- external_connection.export
		);

	mult : component MySoc_m
		port map (
			clk        => clk_clk,                                                --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mult_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => mult_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => mult_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => mult_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => mult_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => mult_export                                             -- external_connection.export
		);

	res : component MySoc_res
		port map (
			clk      => clk_clk,                                        --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => res_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => res_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => res_export                                      -- external_connection.export
		);

	prt : component MySoc_prt
		port map (
			clk      => clk_clk,                                        --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => prt_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => prt_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => prt_export                                      -- external_connection.export
		);

	go : component MySoc_go
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => go_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => go_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => go_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => go_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => go_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => go_export                                             -- external_connection.export
		);

	performance_counter_0 : component MySoc_performance_counter_0
		port map (
			clk           => clk_clk,                                                                          --           clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,                                     --         reset.reset_n
			address       => performance_counter_0_control_slave_translator_avalon_anti_slave_0_address,       -- control_slave.address
			begintransfer => performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer, --              .begintransfer
			readdata      => performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata,      --              .readdata
			write         => performance_counter_0_control_slave_translator_avalon_anti_slave_0_write,         --              .write
			writedata     => performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata      --              .writedata
		);

	nios_instruction_master_translator : component mysoc_nios_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 18,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 18,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                    --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                             --                     reset.reset
			uav_address              => nios_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => nios_instruction_master_read,                                               --                          .read
			av_readdata              => nios_instruction_master_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                        --               (terminated)
			av_byteenable            => "1111",                                                                     --               (terminated)
			av_beginbursttransfer    => '0',                                                                        --               (terminated)
			av_begintransfer         => '0',                                                                        --               (terminated)
			av_chipselect            => '0',                                                                        --               (terminated)
			av_readdatavalid         => open,                                                                       --               (terminated)
			av_write                 => '0',                                                                        --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                         --               (terminated)
			av_lock                  => '0',                                                                        --               (terminated)
			av_debugaccess           => '0',                                                                        --               (terminated)
			uav_clken                => open,                                                                       --               (terminated)
			av_clken                 => '1',                                                                        --               (terminated)
			uav_response             => "00",                                                                       --               (terminated)
			av_response              => open,                                                                       --               (terminated)
			uav_writeresponserequest => open,                                                                       --               (terminated)
			uav_writeresponsevalid   => '0',                                                                        --               (terminated)
			av_writeresponserequest  => '0',                                                                        --               (terminated)
			av_writeresponsevalid    => open                                                                        --               (terminated)
		);

	nios_data_master_translator : component mysoc_nios_data_master_translator
		generic map (
			AV_ADDRESS_W                => 18,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 18,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => clk_clk,                                                             --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                     reset.reset
			uav_address              => nios_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => nios_data_master_byteenable,                                         --                          .byteenable
			av_read                  => nios_data_master_read,                                               --                          .read
			av_readdata              => nios_data_master_readdata,                                           --                          .readdata
			av_write                 => nios_data_master_write,                                              --                          .write
			av_writedata             => nios_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => nios_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                 --               (terminated)
			av_beginbursttransfer    => '0',                                                                 --               (terminated)
			av_begintransfer         => '0',                                                                 --               (terminated)
			av_chipselect            => '0',                                                                 --               (terminated)
			av_readdatavalid         => open,                                                                --               (terminated)
			av_lock                  => '0',                                                                 --               (terminated)
			uav_clken                => open,                                                                --               (terminated)
			av_clken                 => '1',                                                                 --               (terminated)
			uav_response             => "00",                                                                --               (terminated)
			av_response              => open,                                                                --               (terminated)
			uav_writeresponserequest => open,                                                                --               (terminated)
			uav_writeresponsevalid   => '0',                                                                 --               (terminated)
			av_writeresponserequest  => '0',                                                                 --               (terminated)
			av_writeresponsevalid    => open                                                                 --               (terminated)
		);

	nios_jtag_debug_module_translator : component mysoc_nios_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                    --                    reset.reset
			uav_address              => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => nios_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => nios_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => nios_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => nios_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => nios_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => nios_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => nios_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => nios_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_readdatavalid         => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			av_chipselect            => open,                                                                              --              (terminated)
			av_clken                 => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	ram_s1_translator : component mysoc_ram_s1_translator
		generic map (
			AV_ADDRESS_W                   => 14,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                --                    reset.reset
			uav_address              => ram_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ram_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ram_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ram_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ram_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => ram_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => ram_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => ram_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => ram_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => ram_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => ram_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                              --              (terminated)
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	jtag_avalon_jtag_slave_translator : component mysoc_jtag_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                --                    reset.reset
			uav_address              => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_byteenable            => open,                                                                              --              (terminated)
			av_readdatavalid         => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			av_clken                 => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_debugaccess           => open,                                                                              --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	sysid_control_slave_translator : component mysoc_sysid_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                             --                    reset.reset
			uav_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                           --              (terminated)
			av_read                  => open,                                                                           --              (terminated)
			av_writedata             => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	performance_counter_0_control_slave_translator : component mysoc_performance_counter_0_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                        --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                             --                    reset.reset
			uav_address              => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => performance_counter_0_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => performance_counter_0_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_read                  => open,                                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                                           --              (terminated)
			av_burstcount            => open,                                                                                           --              (terminated)
			av_byteenable            => open,                                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                                           --              (terminated)
			av_lock                  => open,                                                                                           --              (terminated)
			av_chipselect            => open,                                                                                           --              (terminated)
			av_clken                 => open,                                                                                           --              (terminated)
			uav_clken                => '0',                                                                                            --              (terminated)
			av_debugaccess           => open,                                                                                           --              (terminated)
			av_outputenable          => open,                                                                                           --              (terminated)
			uav_response             => open,                                                                                           --              (terminated)
			av_response              => "00",                                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                                             --              (terminated)
		);

	m_s1_translator : component mysoc_m_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                         --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                              --                    reset.reset
			uav_address              => m_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => m_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => m_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => m_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => m_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => m_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => m_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => m_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => m_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => m_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => m_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => m_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => m_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => m_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => m_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => m_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                            --              (terminated)
			av_begintransfer         => open,                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                            --              (terminated)
			av_burstcount            => open,                                                            --              (terminated)
			av_byteenable            => open,                                                            --              (terminated)
			av_readdatavalid         => '0',                                                             --              (terminated)
			av_waitrequest           => '0',                                                             --              (terminated)
			av_writebyteenable       => open,                                                            --              (terminated)
			av_lock                  => open,                                                            --              (terminated)
			av_clken                 => open,                                                            --              (terminated)
			uav_clken                => '0',                                                             --              (terminated)
			av_debugaccess           => open,                                                            --              (terminated)
			av_outputenable          => open,                                                            --              (terminated)
			uav_response             => open,                                                            --              (terminated)
			av_response              => "00",                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                            --              (terminated)
			av_writeresponserequest  => open,                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                              --              (terminated)
		);

	mult_s1_translator : component mysoc_m_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                            --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                 --                    reset.reset
			uav_address              => mult_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => mult_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => mult_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => mult_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => mult_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => mult_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => mult_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => mult_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => mult_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => mult_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => mult_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => mult_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => mult_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => mult_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => mult_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => mult_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                               --              (terminated)
			av_begintransfer         => open,                                                               --              (terminated)
			av_beginbursttransfer    => open,                                                               --              (terminated)
			av_burstcount            => open,                                                               --              (terminated)
			av_byteenable            => open,                                                               --              (terminated)
			av_readdatavalid         => '0',                                                                --              (terminated)
			av_waitrequest           => '0',                                                                --              (terminated)
			av_writebyteenable       => open,                                                               --              (terminated)
			av_lock                  => open,                                                               --              (terminated)
			av_clken                 => open,                                                               --              (terminated)
			uav_clken                => '0',                                                                --              (terminated)
			av_debugaccess           => open,                                                               --              (terminated)
			av_outputenable          => open,                                                               --              (terminated)
			uav_response             => open,                                                               --              (terminated)
			av_response              => "00",                                                               --              (terminated)
			uav_writeresponserequest => '0',                                                                --              (terminated)
			uav_writeresponsevalid   => open,                                                               --              (terminated)
			av_writeresponserequest  => open,                                                               --              (terminated)
			av_writeresponsevalid    => '0'                                                                 --              (terminated)
		);

	res_s1_translator : component mysoc_res_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                --                    reset.reset
			uav_address              => res_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => res_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => res_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => res_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => res_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => res_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => res_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => res_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => res_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => res_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => res_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => res_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => res_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                              --              (terminated)
			av_read                  => open,                                                              --              (terminated)
			av_writedata             => open,                                                              --              (terminated)
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_chipselect            => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	prt_s1_translator : component mysoc_res_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                --                    reset.reset
			uav_address              => prt_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => prt_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => prt_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => prt_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => prt_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => prt_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => prt_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => prt_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => prt_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => prt_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => prt_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => prt_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => prt_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                              --              (terminated)
			av_read                  => open,                                                              --              (terminated)
			av_writedata             => open,                                                              --              (terminated)
			av_begintransfer         => open,                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_chipselect            => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	go_s1_translator : component mysoc_m_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 18,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                          --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                               --                    reset.reset
			uav_address              => go_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => go_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => go_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => go_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => go_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => go_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => go_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => go_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => go_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => go_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => go_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => go_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => go_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => go_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => go_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => go_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                             --              (terminated)
			av_begintransfer         => open,                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                             --              (terminated)
			av_burstcount            => open,                                                             --              (terminated)
			av_byteenable            => open,                                                             --              (terminated)
			av_readdatavalid         => '0',                                                              --              (terminated)
			av_waitrequest           => '0',                                                              --              (terminated)
			av_writebyteenable       => open,                                                             --              (terminated)
			av_lock                  => open,                                                             --              (terminated)
			av_clken                 => open,                                                             --              (terminated)
			uav_clken                => '0',                                                              --              (terminated)
			av_debugaccess           => open,                                                             --              (terminated)
			av_outputenable          => open,                                                             --              (terminated)
			uav_response             => open,                                                             --              (terminated)
			av_response              => "00",                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                             --              (terminated)
			av_writeresponserequest  => open,                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                               --              (terminated)
		);

	nios_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_BEGIN_BURST           => 73,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			PKT_BURST_TYPE_H          => 70,
			PKT_BURST_TYPE_L          => 69,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_TRANS_EXCLUSIVE       => 59,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_THREAD_ID_H           => 83,
			PKT_THREAD_ID_L           => 83,
			PKT_CACHE_H               => 90,
			PKT_CACHE_L               => 87,
			PKT_DATA_SIDEBAND_H       => 72,
			PKT_DATA_SIDEBAND_L       => 72,
			PKT_QOS_H                 => 74,
			PKT_QOS_L                 => 74,
			PKT_ADDR_SIDEBAND_H       => 71,
			PKT_ADDR_SIDEBAND_L       => 71,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			ST_DATA_W                 => 93,
			ST_CHANNEL_W              => 10,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                             --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			av_address              => nios_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                              --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                               --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                            --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                      --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                        --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                              --          .ready
			av_response             => open,                                                                                -- (terminated)
			av_writeresponserequest => '0',                                                                                 -- (terminated)
			av_writeresponsevalid   => open                                                                                 -- (terminated)
		);

	nios_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_BEGIN_BURST           => 73,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			PKT_BURST_TYPE_H          => 70,
			PKT_BURST_TYPE_L          => 69,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_TRANS_EXCLUSIVE       => 59,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_THREAD_ID_H           => 83,
			PKT_THREAD_ID_L           => 83,
			PKT_CACHE_H               => 90,
			PKT_CACHE_L               => 87,
			PKT_DATA_SIDEBAND_H       => 72,
			PKT_DATA_SIDEBAND_L       => 72,
			PKT_QOS_H                 => 74,
			PKT_QOS_L                 => 74,
			PKT_ADDR_SIDEBAND_H       => 71,
			PKT_ADDR_SIDEBAND_L       => 71,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			ST_DATA_W                 => 93,
			ST_CHANNEL_W              => 10,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                      --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			av_address              => nios_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                   --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                    --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                 --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                           --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                             --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                   --          .ready
			av_response             => open,                                                                         -- (terminated)
			av_writeresponserequest => '0',                                                                          -- (terminated)
			av_writeresponsevalid   => open                                                                          -- (terminated)
		);

	nios_jtag_debug_module_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                              --       clk_reset.reset
			m0_address              => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                      --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                    --                .channel
			rf_sink_ready           => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                          --     (terminated)
		);

	nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			in_data           => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	ram_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                          --       clk_reset.reset
			m0_address              => ram_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ram_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ram_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ram_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ram_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ram_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ram_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                --                .channel
			rf_sink_ready           => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			in_data           => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_002_src_ready,                                                                  --              cp.ready
			cp_valid                => cmd_xbar_mux_002_src_valid,                                                                  --                .valid
			cp_data                 => cmd_xbar_mux_002_src_data,                                                                   --                .data
			cp_startofpacket        => cmd_xbar_mux_002_src_startofpacket,                                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_002_src_endofpacket,                                                            --                .endofpacket
			cp_channel              => cmd_xbar_mux_002_src_channel,                                                                --                .channel
			rf_sink_ready           => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                          --     (terminated)
		);

	jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                       --       clk_reset.reset
			m0_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_003_src_ready,                                                               --              cp.ready
			cp_valid                => cmd_xbar_mux_003_src_valid,                                                               --                .valid
			cp_data                 => cmd_xbar_mux_003_src_data,                                                                --                .data
			cp_startofpacket        => cmd_xbar_mux_003_src_startofpacket,                                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_003_src_endofpacket,                                                         --                .endofpacket
			cp_channel              => cmd_xbar_mux_003_src_channel,                                                             --                .channel
			rf_sink_ready           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                  --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                                  --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                       --       clk_reset.reset
			m0_address              => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_004_src_ready,                                                                               --              cp.ready
			cp_valid                => cmd_xbar_mux_004_src_valid,                                                                               --                .valid
			cp_data                 => cmd_xbar_mux_004_src_data,                                                                                --                .data
			cp_startofpacket        => cmd_xbar_mux_004_src_startofpacket,                                                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_004_src_endofpacket,                                                                         --                .endofpacket
			cp_channel              => cmd_xbar_mux_004_src_channel,                                                                             --                .channel
			rf_sink_ready           => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                       --     (terminated)
		);

	performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                                  --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                       -- clk_reset.reset
			in_data           => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                     -- (terminated)
			csr_read          => '0',                                                                                                      -- (terminated)
			csr_write         => '0',                                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                       -- (terminated)
			almost_full_data  => open,                                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                                     -- (terminated)
			in_empty          => '0',                                                                                                      -- (terminated)
			out_empty         => open,                                                                                                     -- (terminated)
			in_error          => '0',                                                                                                      -- (terminated)
			out_error         => open,                                                                                                     -- (terminated)
			in_channel        => '0',                                                                                                      -- (terminated)
			out_channel       => open                                                                                                      -- (terminated)
		);

	m_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                   --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                        --       clk_reset.reset
			m0_address              => m_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => m_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => m_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => m_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => m_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => m_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => m_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => m_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => m_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => m_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => m_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => m_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => m_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => m_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => m_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => m_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src5_ready,                                             --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src5_valid,                                             --                .valid
			cp_data                 => cmd_xbar_demux_001_src5_data,                                              --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src5_startofpacket,                                     --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src5_endofpacket,                                       --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src5_channel,                                           --                .channel
			rf_sink_ready           => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => m_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => m_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => m_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => m_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => m_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => m_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                        --     (terminated)
		);

	m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                   --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                        -- clk_reset.reset
			in_data           => m_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => m_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => m_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => m_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => m_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => m_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                      -- (terminated)
			csr_read          => '0',                                                                       -- (terminated)
			csr_write         => '0',                                                                       -- (terminated)
			csr_readdata      => open,                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                        -- (terminated)
			almost_full_data  => open,                                                                      -- (terminated)
			almost_empty_data => open,                                                                      -- (terminated)
			in_empty          => '0',                                                                       -- (terminated)
			out_empty         => open,                                                                      -- (terminated)
			in_error          => '0',                                                                       -- (terminated)
			out_error         => open,                                                                      -- (terminated)
			in_channel        => '0',                                                                       -- (terminated)
			out_channel       => open                                                                       -- (terminated)
		);

	mult_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                           --       clk_reset.reset
			m0_address              => mult_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => mult_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => mult_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => mult_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => mult_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => mult_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => mult_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => mult_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => mult_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => mult_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => mult_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => mult_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => mult_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => mult_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => mult_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => mult_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src6_ready,                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src6_valid,                                                --                .valid
			cp_data                 => cmd_xbar_demux_001_src6_data,                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src6_startofpacket,                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src6_endofpacket,                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src6_channel,                                              --                .channel
			rf_sink_ready           => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => mult_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                         --     (terminated)
			m0_writeresponserequest => open,                                                                         --     (terminated)
			m0_writeresponsevalid   => '0'                                                                           --     (terminated)
		);

	mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                           -- clk_reset.reset
			in_data           => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => mult_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => mult_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                         -- (terminated)
			csr_read          => '0',                                                                          -- (terminated)
			csr_write         => '0',                                                                          -- (terminated)
			csr_readdata      => open,                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                           -- (terminated)
			almost_full_data  => open,                                                                         -- (terminated)
			almost_empty_data => open,                                                                         -- (terminated)
			in_empty          => '0',                                                                          -- (terminated)
			out_empty         => open,                                                                         -- (terminated)
			in_error          => '0',                                                                          -- (terminated)
			out_error         => open,                                                                         -- (terminated)
			in_channel        => '0',                                                                          -- (terminated)
			out_channel       => open                                                                          -- (terminated)
		);

	res_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                          --       clk_reset.reset
			m0_address              => res_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => res_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => res_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => res_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => res_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => res_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => res_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => res_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => res_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => res_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => res_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => res_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => res_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => res_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => res_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => res_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                               --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                               --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                                --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                         --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                             --                .channel
			rf_sink_ready           => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => res_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => res_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => res_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => res_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => res_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => res_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			in_data           => res_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => res_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => res_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => res_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => res_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => res_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	prt_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                          --       clk_reset.reset
			m0_address              => prt_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => prt_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => prt_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => prt_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => prt_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => prt_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => prt_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => prt_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => prt_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => prt_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => prt_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => prt_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => prt_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => prt_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => prt_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => prt_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src8_ready,                                               --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src8_valid,                                               --                .valid
			cp_data                 => cmd_xbar_demux_001_src8_data,                                                --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src8_startofpacket,                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src8_endofpacket,                                         --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src8_channel,                                             --                .channel
			rf_sink_ready           => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => prt_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                          --     (terminated)
		);

	prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                          -- clk_reset.reset
			in_data           => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => prt_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => prt_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                        -- (terminated)
			csr_read          => '0',                                                                         -- (terminated)
			csr_write         => '0',                                                                         -- (terminated)
			csr_readdata      => open,                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                          -- (terminated)
			almost_full_data  => open,                                                                        -- (terminated)
			almost_empty_data => open,                                                                        -- (terminated)
			in_empty          => '0',                                                                         -- (terminated)
			out_empty         => open,                                                                        -- (terminated)
			in_error          => '0',                                                                         -- (terminated)
			out_error         => open,                                                                        -- (terminated)
			in_channel        => '0',                                                                         -- (terminated)
			out_channel       => open                                                                         -- (terminated)
		);

	go_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 73,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 53,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 54,
			PKT_TRANS_POSTED          => 55,
			PKT_TRANS_WRITE           => 56,
			PKT_TRANS_READ            => 57,
			PKT_TRANS_LOCK            => 58,
			PKT_SRC_ID_H              => 78,
			PKT_SRC_ID_L              => 75,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 79,
			PKT_BURSTWRAP_H           => 65,
			PKT_BURSTWRAP_L           => 63,
			PKT_BYTE_CNT_H            => 62,
			PKT_BYTE_CNT_L            => 60,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 68,
			PKT_BURST_SIZE_L          => 66,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                    --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                         --       clk_reset.reset
			m0_address              => go_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => go_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => go_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => go_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => go_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => go_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => go_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => go_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => go_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => go_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => go_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => go_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => go_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => go_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => go_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => go_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src9_ready,                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src9_valid,                                              --                .valid
			cp_data                 => cmd_xbar_demux_001_src9_data,                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src9_startofpacket,                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src9_endofpacket,                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src9_channel,                                            --                .channel
			rf_sink_ready           => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => go_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => go_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => go_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => go_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => go_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => go_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                         --     (terminated)
		);

	go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 94,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                         -- clk_reset.reset
			in_data           => go_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => go_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => go_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => go_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => go_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => go_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                       -- (terminated)
			csr_read          => '0',                                                                        -- (terminated)
			csr_write         => '0',                                                                        -- (terminated)
			csr_readdata      => open,                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                         -- (terminated)
			almost_full_data  => open,                                                                       -- (terminated)
			almost_empty_data => open,                                                                       -- (terminated)
			in_empty          => '0',                                                                        -- (terminated)
			out_empty         => open,                                                                       -- (terminated)
			in_error          => '0',                                                                        -- (terminated)
			out_error         => open,                                                                       -- (terminated)
			in_channel        => '0',                                                                        -- (terminated)
			out_channel       => open                                                                        -- (terminated)
		);

	addr_router : component MySoc_addr_router
		port map (
			sink_ready         => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                               --       src.ready
			src_valid          => addr_router_src_valid,                                                               --          .valid
			src_data           => addr_router_src_data,                                                                --          .data
			src_channel        => addr_router_src_channel,                                                             --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                          --          .endofpacket
		);

	addr_router_001 : component MySoc_addr_router_001
		port map (
			sink_ready         => nios_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                    --       src.ready
			src_valid          => addr_router_001_src_valid,                                                    --          .valid
			src_data           => addr_router_001_src_data,                                                     --          .data
			src_channel        => addr_router_001_src_channel,                                                  --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                            --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                               --          .endofpacket
		);

	id_router : component MySoc_id_router
		port map (
			sink_ready         => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                               --       src.ready
			src_valid          => id_router_src_valid,                                                               --          .valid
			src_data           => id_router_src_data,                                                                --          .data
			src_channel        => id_router_src_channel,                                                             --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                          --          .endofpacket
		);

	id_router_001 : component MySoc_id_router
		port map (
			sink_ready         => ram_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ram_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ram_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                           --       src.ready
			src_valid          => id_router_001_src_valid,                                           --          .valid
			src_data           => id_router_001_src_data,                                            --          .data
			src_channel        => id_router_001_src_channel,                                         --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                      --          .endofpacket
		);

	id_router_002 : component MySoc_id_router
		port map (
			sink_ready         => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                           --       src.ready
			src_valid          => id_router_002_src_valid,                                                           --          .valid
			src_data           => id_router_002_src_data,                                                            --          .data
			src_channel        => id_router_002_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                      --          .endofpacket
		);

	id_router_003 : component MySoc_id_router
		port map (
			sink_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                        --       src.ready
			src_valid          => id_router_003_src_valid,                                                        --          .valid
			src_data           => id_router_003_src_data,                                                         --          .data
			src_channel        => id_router_003_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                   --          .endofpacket
		);

	id_router_004 : component MySoc_id_router
		port map (
			sink_ready         => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                             -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                                        --       src.ready
			src_valid          => id_router_004_src_valid,                                                                        --          .valid
			src_data           => id_router_004_src_data,                                                                         --          .data
			src_channel        => id_router_004_src_channel,                                                                      --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                                --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                                   --          .endofpacket
		);

	id_router_005 : component MySoc_id_router_005
		port map (
			sink_ready         => m_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => m_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => m_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => m_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => m_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                         --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                              -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                         --       src.ready
			src_valid          => id_router_005_src_valid,                                         --          .valid
			src_data           => id_router_005_src_data,                                          --          .data
			src_channel        => id_router_005_src_channel,                                       --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                 --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                    --          .endofpacket
		);

	id_router_006 : component MySoc_id_router_005
		port map (
			sink_ready         => mult_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => mult_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => mult_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => mult_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => mult_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                            --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                 -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                            --       src.ready
			src_valid          => id_router_006_src_valid,                                            --          .valid
			src_data           => id_router_006_src_data,                                             --          .data
			src_channel        => id_router_006_src_channel,                                          --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                    --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                       --          .endofpacket
		);

	id_router_007 : component MySoc_id_router_005
		port map (
			sink_ready         => res_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => res_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => res_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => res_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => res_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                           --       src.ready
			src_valid          => id_router_007_src_valid,                                           --          .valid
			src_data           => id_router_007_src_data,                                            --          .data
			src_channel        => id_router_007_src_channel,                                         --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                      --          .endofpacket
		);

	id_router_008 : component MySoc_id_router_005
		port map (
			sink_ready         => prt_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => prt_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => prt_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => prt_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => prt_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                           --       src.ready
			src_valid          => id_router_008_src_valid,                                           --          .valid
			src_data           => id_router_008_src_data,                                            --          .data
			src_channel        => id_router_008_src_channel,                                         --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                   --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                      --          .endofpacket
		);

	id_router_009 : component MySoc_id_router_005
		port map (
			sink_ready         => go_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => go_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => go_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => go_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => go_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                          --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                               -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                          --       src.ready
			src_valid          => id_router_009_src_valid,                                          --          .valid
			src_data           => id_router_009_src_data,                                           --          .data
			src_channel        => id_router_009_src_channel,                                        --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                  --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                     --          .endofpacket
		);

	rst_controller : component mysoc_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component mysoc_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1  => nios_jtag_debug_module_reset_reset,     -- reset_in1.reset
			clk        => clk_clk,                                --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req  => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_in2  => '0',                                    -- (terminated)
			reset_in3  => '0',                                    -- (terminated)
			reset_in4  => '0',                                    -- (terminated)
			reset_in5  => '0',                                    -- (terminated)
			reset_in6  => '0',                                    -- (terminated)
			reset_in7  => '0',                                    -- (terminated)
			reset_in8  => '0',                                    -- (terminated)
			reset_in9  => '0',                                    -- (terminated)
			reset_in10 => '0',                                    -- (terminated)
			reset_in11 => '0',                                    -- (terminated)
			reset_in12 => '0',                                    -- (terminated)
			reset_in13 => '0',                                    -- (terminated)
			reset_in14 => '0',                                    -- (terminated)
			reset_in15 => '0'                                     -- (terminated)
		);

	cmd_xbar_demux : component MySoc_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket,   --          .endofpacket
			src3_ready         => cmd_xbar_demux_src3_ready,         --      src3.ready
			src3_valid         => cmd_xbar_demux_src3_valid,         --          .valid
			src3_data          => cmd_xbar_demux_src3_data,          --          .data
			src3_channel       => cmd_xbar_demux_src3_channel,       --          .channel
			src3_startofpacket => cmd_xbar_demux_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_src3_endofpacket,   --          .endofpacket
			src4_ready         => cmd_xbar_demux_src4_ready,         --      src4.ready
			src4_valid         => cmd_xbar_demux_src4_valid,         --          .valid
			src4_data          => cmd_xbar_demux_src4_data,          --          .data
			src4_channel       => cmd_xbar_demux_src4_channel,       --          .channel
			src4_startofpacket => cmd_xbar_demux_src4_startofpacket, --          .startofpacket
			src4_endofpacket   => cmd_xbar_demux_src4_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component MySoc_cmd_xbar_demux_001
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_001_src_ready,             --      sink.ready
			sink_channel       => addr_router_001_src_channel,           --          .channel
			sink_data          => addr_router_001_src_data,              --          .data
			sink_startofpacket => addr_router_001_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_001_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_001_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket,   --          .endofpacket
			src3_ready         => cmd_xbar_demux_001_src3_ready,         --      src3.ready
			src3_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			src3_data          => cmd_xbar_demux_001_src3_data,          --          .data
			src3_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			src3_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_001_src3_endofpacket,   --          .endofpacket
			src4_ready         => cmd_xbar_demux_001_src4_ready,         --      src4.ready
			src4_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			src4_data          => cmd_xbar_demux_001_src4_data,          --          .data
			src4_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			src4_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			src4_endofpacket   => cmd_xbar_demux_001_src4_endofpacket,   --          .endofpacket
			src5_ready         => cmd_xbar_demux_001_src5_ready,         --      src5.ready
			src5_valid         => cmd_xbar_demux_001_src5_valid,         --          .valid
			src5_data          => cmd_xbar_demux_001_src5_data,          --          .data
			src5_channel       => cmd_xbar_demux_001_src5_channel,       --          .channel
			src5_startofpacket => cmd_xbar_demux_001_src5_startofpacket, --          .startofpacket
			src5_endofpacket   => cmd_xbar_demux_001_src5_endofpacket,   --          .endofpacket
			src6_ready         => cmd_xbar_demux_001_src6_ready,         --      src6.ready
			src6_valid         => cmd_xbar_demux_001_src6_valid,         --          .valid
			src6_data          => cmd_xbar_demux_001_src6_data,          --          .data
			src6_channel       => cmd_xbar_demux_001_src6_channel,       --          .channel
			src6_startofpacket => cmd_xbar_demux_001_src6_startofpacket, --          .startofpacket
			src6_endofpacket   => cmd_xbar_demux_001_src6_endofpacket,   --          .endofpacket
			src7_ready         => cmd_xbar_demux_001_src7_ready,         --      src7.ready
			src7_valid         => cmd_xbar_demux_001_src7_valid,         --          .valid
			src7_data          => cmd_xbar_demux_001_src7_data,          --          .data
			src7_channel       => cmd_xbar_demux_001_src7_channel,       --          .channel
			src7_startofpacket => cmd_xbar_demux_001_src7_startofpacket, --          .startofpacket
			src7_endofpacket   => cmd_xbar_demux_001_src7_endofpacket,   --          .endofpacket
			src8_ready         => cmd_xbar_demux_001_src8_ready,         --      src8.ready
			src8_valid         => cmd_xbar_demux_001_src8_valid,         --          .valid
			src8_data          => cmd_xbar_demux_001_src8_data,          --          .data
			src8_channel       => cmd_xbar_demux_001_src8_channel,       --          .channel
			src8_startofpacket => cmd_xbar_demux_001_src8_startofpacket, --          .startofpacket
			src8_endofpacket   => cmd_xbar_demux_001_src8_endofpacket,   --          .endofpacket
			src9_ready         => cmd_xbar_demux_001_src9_ready,         --      src9.ready
			src9_valid         => cmd_xbar_demux_001_src9_valid,         --          .valid
			src9_data          => cmd_xbar_demux_001_src9_data,          --          .data
			src9_channel       => cmd_xbar_demux_001_src9_channel,       --          .channel
			src9_startofpacket => cmd_xbar_demux_001_src9_startofpacket, --          .startofpacket
			src9_endofpacket   => cmd_xbar_demux_001_src9_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component MySoc_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component MySoc_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component MySoc_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src2_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src2_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src2_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src2_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src2_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src2_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component MySoc_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_003_src_data,             --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src3_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src3_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src3_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src3_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src3_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src3_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src3_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src3_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_004 : component MySoc_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_004_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_004_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_004_src_data,             --          .data
			src_channel         => cmd_xbar_mux_004_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_004_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_004_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src4_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src4_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src4_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src4_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src4_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src4_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src4_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src4_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src4_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component MySoc_rsp_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component MySoc_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component MySoc_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component MySoc_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component MySoc_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_004_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_004_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_004_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component MySoc_rsp_xbar_demux_005
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component MySoc_rsp_xbar_demux_005
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component MySoc_rsp_xbar_demux_005
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component MySoc_rsp_xbar_demux_005
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component MySoc_rsp_xbar_demux_005
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component MySoc_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component MySoc_rsp_xbar_mux_001
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src1_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src1_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src1_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src1_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src1_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src1_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src1_endofpacket,   --          .endofpacket
			sink5_ready         => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data          => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready         => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready         => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data          => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket   => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready         => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data          => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket   => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready         => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data          => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	irq_mapper : component MySoc_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios_d_irq_irq                  --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	m_s1_translator_avalon_anti_slave_0_write_ports_inv <= not m_s1_translator_avalon_anti_slave_0_write;

	mult_s1_translator_avalon_anti_slave_0_write_ports_inv <= not mult_s1_translator_avalon_anti_slave_0_write;

	go_s1_translator_avalon_anti_slave_0_write_ports_inv <= not go_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of MySoc
