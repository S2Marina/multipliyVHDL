library verilog;
use verilog.vl_types.all;
entity MySoc_nios_nios2_performance_monitors is
end MySoc_nios_nios2_performance_monitors;
